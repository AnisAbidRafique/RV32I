`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/25/2024 11:50:06 PM
// Design Name: 
// Module Name: data_mem_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module data_mem_tb;

    logic [32 - 1 : 0] addr;
    logic [32 - 1 : 0]dataW;
    logic MemRW;
    logic clk;
    logic [2:0] funct3;
    logic [32 - 1 : 0]dataR;

data_mem #(.IMEM_DEPTH(),.PROG_VALUE())  
uutgen
(   .addr(addr),
    .dataW(dataW),
    .MemRW(MemRW),
    .clk(clk),
    .funct3(funct3),
    .dataR(dataR)
);

always #5 clk = ~clk;

// Test bench
initial 
begin
    clk = 0;
    MemRW = 0;
    #10
    
    
    //load byte cases
    funct3 = 0;
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    //addr = 1;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    // addr = 5;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
    // addr = 10;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    // addr = 14;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    // addr = 17;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
    // addr = 22;  
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
    // addr = 25;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0010;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0011;
    
    //load byte unsigned
    #10
    funct3 = 4;
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    //addr = 1;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    // addr = 5;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
    // addr = 10;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    // addr = 14;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    // addr = 17;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
    // addr = 22;  
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
    // addr = 25;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0010;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0011;
    
    //load half byte
    #10
    funct3 = 1;
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    //addr = 1;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    // addr = 5;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
    // addr = 10;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    // addr = 14;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    // addr = 17;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
    // addr = 22;  
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
    // addr = 25;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0010;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0011;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0111;

    //load half byte unsigned
    #10
    funct3 = 5;
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    //addr = 1;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    // addr = 5;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
    // addr = 10;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    // addr = 14;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    // addr = 17;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
    // addr = 22;  
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
    // addr = 25;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0010;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0011;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0111;

    //store instructions
    //store word
    #10
    MemRW = 1;
    funct3 = 2;
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    dataW = 32'hEDCF_1254;
    addr = 1;
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    dataW = 32'hEDCF_0054;
    addr = 5;
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
    dataW = 32'h0DCF_1254;
    addr = 10;
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    dataW = 32'hEDC1_1254;
    addr = 14;
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    dataW = 32'hEDCF_1554;
    addr = 17;
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
    dataW = 32'h7DCF_1254;
    addr = 22;  
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
    dataW = 32'h4DCF_1254;
    addr = 25;
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0010;
    dataW = 32'hEDCF_1274;
    addr = 31;
    #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0011;
    dataW = 32'hEDCF_1284;
    addr = 33;

    #10 
    MemRW = 0;
    addr = 36;

    // //store byte
    // #10
    // funct3 = 0;
    // MemRW  = 1;
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    // dataW = 32'hEDCF_1254;
    // //addr = 1;
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    // dataW = 32'hEDCF_1254;
    // // addr = 5;
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
    // dataW = 32'hEDCF_1254;
    // // addr = 10;
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    // dataW = 32'hEDCF_1254;
    // // addr = 14;
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    // dataW = 32'hEDCF_1254;
    // // addr = 17;
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
    // dataW = 32'hEDCF_1254;
    // // addr = 22;  
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
    // dataW = 32'hEDCF_1254;
    // // addr = 25;
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0010;
    // dataW = 32'hEDCF_1254;
    // #10
    // addr = 32'b0000_0000_0000_0000_0000_0000_0001_0011;
    // dataW = 32'hEDCF_1254;

    //store half byte
    #10
    MemRW  = 1;
    funct3 = 1;
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0001;
    dataW = 32'hEDCF_1254;
    //addr = 1;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0110;
    dataW = 32'hEDCF_1254;
    // addr = 5;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
    dataW = 32'hEDCF_1254;
    // addr = 10;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
    dataW = 32'hEDCF_1254;
    // addr = 14;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0000_0010;
    dataW = 32'hEDCF_1254;
    // addr = 17;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0000;
    dataW = 32'hEDCF_1254;
    // addr = 22;  
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0001;
    dataW = 32'hEDCF_1254;
    // addr = 25;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0010;
    dataW = 32'hEDCF_1254;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0011;
    dataW = 32'hEDCF_1254;
    #10
    addr = 32'b0000_0000_0000_0000_0000_0000_0001_0111;
    dataW = 32'hEDCF_1254;

    #10 
        $stop;
end
endmodule
